 `define DELAY 20
module _32bit_testbench(); 
reg [31:0] a,b;
reg [2:0] op;
wire [31:0] sum;

elveda g1(a,b,op,sum);
initial begin
a = 32'b00000000000000000000000000000011; b = 32'b00000000000000000000000000000001; op = 000;
#`DELAY;
a = 32'b11111000000000000000000000000011; b = 32'b11111111111111111111111111111111; op = 001;
#`DELAY;
a = 32'b00000000000000000000000000000011; b = 32'b00000000000000000000000000000001; op = 010;
#`DELAY;
a = 32'b00000000000000000000000000000000; b = 32'b00000000000000000000000000000001; op = 100;
#`DELAY;
a = 32'b10000000000000000000000000000000; b = 32'b00000000000000000000000000000001; op = 100;
#`DELAY;
a = 32'b10010101000000000000000000000000; b = 32'b11111100101000000000000000000001; op = 101;
#`DELAY;
a = 32'b10010101000000000000000000000000; b = 32'b11111100101000000000000000000001; op = 110;
#`DELAY;
a = 32'b10010101000000000000000000000000; b = 32'b11111100101000000000000000000001; op = 111;
#`DELAY;
end
 
 
initial
begin
$monitor("time = %2d, a =%32b, b=%32b, op=%3b, sum=%32b", $time, a, b, op, sum);
end
 
endmodule
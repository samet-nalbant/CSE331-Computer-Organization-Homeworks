module to32bit_zeros(D,B);
input D;
output [31:0] B;

	or g31(B[31],0,0);
	or g30(B[30],0,0);
	or g29(B[29],0,0);	
	or g28(B[28],0,0);
	
	or g27(B[27],0,0);
	or g26(B[26],0,0);
	or g25(B[25],0,0);	
	or g24(B[24],0,0);
	
	or g23(B[23],0,0);
	or g22(B[22],0,0);
	or g21(B[21],0,0);	
	or g20(B[20],0,0);
	
	or g19(B[19],0,0);
	or g18(B[18],0,0);
	or g17(B[17],0,0);	
	or g16(B[16],0,0);
	
	or g15(B[15],0,0);
	or g14(B[14],0,0);
	or g13(B[13],0,0);	
	or g12(B[12],0,0);
	
	or g11(B[11],0,0);
	or g10(B[10],0,0);
	or g9(B[9],0,0);	
	or g8(B[8],0,0);

	or g7(B[7],0,0);
	or g6(B[6],0,0);
	or g5(B[5],0,0);	
	or g4(B[4],0,0);
	
	or g3(B[3],0,0);
	or g2(B[2],0,0);
	or g1(B[1],0,0);	
	or g0(B[0],D,0);


endmodule 
`define DELAY 20
module _32bit_slt_testbench(); 
reg [31:0] a,b,c,d,e,f,g,h;
reg [2:0]S;
wire [31:0] sum;

elveda g1(a,b,c,d,e,f,g,h,S,sum);
initial begin
a = 32'b11100000000000000000000000000011; b = 32'b00000000000000000000000000000001;c = 32'b00000000000000000000000000000011; d = 32'b00000000000000000000000000000001; e = 32'b00000000000000000000000000000011; f = 32'b00000000000000000000000000000001; g = 32'b00000000000000000000000000000011; h = 32'b00000000000000000000000000000001; S = 000; 
#`DELAY;
a = 32'b00000000000000000000000000000011; b = 32'b10100000000000000000000000000001;c = 32'b00000000000000000000000000000011; d = 32'b00000000000000000000000000000001; e = 32'b00000000000000000000000000000011; f = 32'b00000000000000000000000000000001; g = 32'b00000000000000000000000000000011; h = 32'b00000000000000000000000000000001; S = 001;
#`DELAY;
end
 
 
initial
begin
$monitor("time = %2d, sum=%32b", $time,sum);
end
 
endmodule